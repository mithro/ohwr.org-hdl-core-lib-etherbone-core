---! Standard library
library IEEE;
--! Standard packages    
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.vhdl_2008_workaround_pkg.all;

entity WB_bus_adapter is
generic(g_adr_width_A : natural := 32; g_adr_width_B  : natural := 32;
		g_dat_width_A : natural := 32; g_dat_width_B  : natural := 16;
		g_pipeline : natural 
		);
		-- pipeline: 0 => A-x, 1 x-B, 2 A-B 
port(
		clk_i		: in std_logic;
		nRst_i		: in std_logic;
		
		A_CYC_i		: in std_logic;
		A_STB_i		: in std_logic;
		A_ADR_i		: in std_logic_vector(g_adr_width_A-1 downto 0);
		A_SEL_i		: in std_logic_vector(g_dat_width_A/8-1 downto 0);
		A_WE_i		: in std_logic;
		A_DAT_i		: in std_logic_vector(g_dat_width_A-1 downto 0);
		A_ACK_o		: out std_logic;
		A_ERR_o		: out std_logic;
		A_RTY_o		: out std_logic;
		A_STALL_o	: out std_logic;
		A_DAT_o		: out std_logic_vector(g_dat_width_A-1 downto 0);
		
		
		B_CYC_o		: out std_logic;
		B_STB_o		: out std_logic;
		B_ADR_o		: out std_logic_vector(g_adr_width_B-1 downto 0);
		B_SEL_o		: out std_logic_vector(g_dat_width_B/8-1 downto 0);
		B_WE_o		: out std_logic;
		B_DAT_o		: out std_logic_vector(g_dat_width_B-1 downto 0);
		B_ACK_i		: in std_logic;
		B_ERR_i		: in std_logic;
		B_RTY_i		: in std_logic;
		B_STALL_i	: in std_logic;
		B_DAT_i		: in std_logic_vector(g_dat_width_B-1 downto 0)

);
end WB_bus_adapter;




architecture behavioral of WB_bus_adapter is

	constant c_adr_w_max : natural := maximum(g_adr_width_A, g_adr_width_B);
	constant c_dat_w_max : natural := maximum(g_dat_width_A, g_dat_width_B);
	constant c_sel_w_max : natural := maximum(g_dat_width_A, g_dat_width_B)/8;
	constant c_adr_w_min : natural := minimum(g_adr_width_A, g_adr_width_B);
	constant c_dat_w_min : natural := minimum(g_dat_width_A, g_dat_width_B);
	constant c_sel_w_min : natural := minimum(g_dat_width_A, g_dat_width_B)/8;
	
	signal sipo_d	 : std_logic_vector(c_dat_w_min-1 downto 0);
	signal sipo_q	 : std_logic_vector(c_dat_w_max-1 downto 0);
	signal piso_d	 : std_logic_vector(c_dat_w_max-1 downto 0);
	signal piso_q	 : std_logic_vector(c_dat_w_min-1 downto 0);
	
	-- direct adapter signals
	constant c_adr_pad 	: std_logic_vector(c_adr_w_max-1 downto 0) 	:=  (others => '0');
	constant c_sel_pad 	: std_logic_vector(c_sel_w_max-1 downto 0) 	:=  (others => '0');
	constant c_dat_pad 	: std_logic_vector(c_dat_w_max-1 downto 0) 	:=  (others => '0');
	
	signal 	adr 		: std_logic_vector(c_adr_w_max-1 downto 0);
	signal 	slave_dat 	: std_logic_vector(c_dat_w_max-1 downto 0);
	signal 	master_dat 	: std_logic_vector(c_dat_w_max-1 downto 0);
	signal 	sel 		: std_logic_vector(c_sel_w_max-1 downto 0);
	signal  cyc : std_logic;
	
	-- S/G adapter signals
	signal sipo_sh_in 	: std_logic;
	signal sipo_clr 	: std_logic;
	signal sipo_full 	: std_logic;
	
	signal piso_sh_out 	: std_logic;
	signal piso_ld 	: std_logic;
	signal piso_empty 	: std_logic;
	signal ld 	: std_logic;
	
	signal get_adr : std_logic;
	
		
	component sipo_flag is
	generic(g_width_IN : natural := 16; g_width_OUT  : natural := 32); 
	port(
			clk_i				: in std_logic;
			nRst_i				: in std_logic;
			
			d_i					: in std_logic_vector(g_width_IN-1 downto 0);
			en_i				: in std_logic;
			clr_i				: in std_logic;
			
			q_o					: out std_logic_vector(g_width_OUT-1 downto 0);
			full_o				: out std_logic

	);
	end component;
	
	component piso_flag is
	generic(g_width_IN : natural := 16; g_width_OUT  : natural := 32); 
	port(
			clk_i				: in std_logic;
			nRst_i				: in std_logic;
			
			d_i					: in std_logic_vector(g_width_IN-1 downto 0);
			en_i				: in std_logic;
			ld_i				: in std_logic;
			
			q_o					: out std_logic_vector(g_width_OUT-1 downto 0);
			empty_o				: out std_logic

	);
	end component;

begin


	
---------------------------------------------------------------------------------------------------------------------------------	
PIPELINED:		if(g_pipeline = 2) GENERATE		
		
		
A_LESSER_B:		if(c_dat_w_min = g_dat_width_A) GENERATE
			gather : sipo_flag -- MA ->-> => MB
			generic map(g_width_IN => c_dat_w_min, g_width_OUT  => c_dat_w_max) 
			port map(
			clk_i		=> clk_i,
			nRst_i	=> nRSt_i,
			
			d_i			=> sipo_d,
			en_i		=> sipo_sh_in,
			clr_i		=> sipo_clr,
			
			q_o			=> sipo_q,
			full_o		=> sipo_full
			);
			
			sipo_d <= A_DAT_i;
			B_DAT_o <= sipo_q;
			B_ADR_o <= adr(B_ADR_o'left downto 0);
			
			scatter : piso_flag -- SB => ->-> SA 
			generic map(g_width_IN => c_dat_w_max, g_width_OUT  => c_dat_w_min) 
			port map(
			clk_i		=> clk_i,
			nRst_i		=> nRSt_i,
			
			d_i			=> piso_d,
			en_i		=> piso_sh_out,
			ld_i		=> piso_ld,
			
			q_o			=> piso_q,
			empty_o		=> piso_empty
			);
		
			-- PISO -- SB => ->-> SA 
			piso_d 		<= B_DAT_i;
			A_DAT_o 	<= piso_q;
			piso_ld 	<= B_ACK_i;
			A_ACK_o 	<= NOT piso_empty;
			piso_sh_out <= NOT piso_empty;
			
			process (clk_i)
			begin
				if (clk_i'event and clk_i = '1') then
					if(nRSt_i = '0') then
						B_CYC_o 	<= '0';
						B_STB_o 	<= '0';
						A_ACK_o 	<= '0';
						A_STALL_o 	<= '0';
						CYC 		<= '0';
						
						piso_ld 	<= '0';
						piso_sh_out	<= '0';
						sipo_clr 	<= '0';
						sipo_sh_in 	<= '0';

					else
						B_CYC_o 	<= '0';
						B_STB_o 	<= '0';
						A_ACK_o 	<= '0';
						A_STALL_o 	<= '0';
						piso_ld 	<= '0';
						piso_sh_out	<= '0';
						sipo_clr 	<= '0';
						sipo_sh_in 	<= '0';
						
						CYC <= A_CYC_i;
						
						-- SIPO -- MA ->-> => MB
						--sipo_clr
						if(sipo_full ='1' AND B_STALL_i = '0') then
							sipo_clr <= '1';
							--get_adr <= '1';
							--adr <= (others => '0');
						end if;	
						
						--adr
						--if(sipo_full ='0' AND get_adr = '1') then
						--	adr(A_ADR_i'left downto ld(g_dat_width_A/8-1)) <= A_ADR_i(A_ADR_i'left downto ld(g_dat_width_A/8-1));
						--	get_adr <= '0'
						--end if;	
						
						--sipo_sh_in
						if(sipo_full ='0') then
							sipo_sh_in <= '1';
						end if;	
						
						-- CYC
						if(A_CYC_i = '1' OR sipo_full= '1') then
							B_CYC_o <= '1';
						end if;
						
						-- STB	
						if((A_CYC_i = '0' AND CYC = '1') OR sipo_full ='1') then--falling edge
							B_STB_o <= '1';
						end if;
						
						-- STALL
						if(sipo_full ='1' AND B_STALL_i = '1') then
							A_STALL_o <= '1';
						end if;	
						
						

						

					end if;	
				end if;
			end process;
				
		END GENERATE;
		
		--scatter
A_GREATER_B:				if(c_dat_w_max = g_dat_width_A) GENERATE
			scatter : piso_flag -- MA => ->-> MB
			generic map(g_width_IN => c_dat_w_max, g_width_OUT  => c_dat_w_min) 
			port map(
			clk_i		=> clk_i,
			nRst_i		=> nRSt_i,
			
			d_i			=> piso_d,
			en_i		=> piso_sh_out,
			ld_i		=> piso_ld,
			
			q_o			=> piso_q,
			empty_o		=> piso_empty
			);
		
			piso_d 		<= A_DAT_i;
			B_DAT_o 	<= piso_q;
			
			
			gather : sipo_flag -- SB ->-> => SA
			generic map(g_width_IN => c_dat_w_min, g_width_OUT  => c_dat_w_max) 
			port map(
			clk_i		=> clk_i,
			nRst_i	=> nRSt_i,
			
			d_i			=> sipo_d,
			en_i		=> sipo_sh_in,
			clr_i		=> sipo_clr,
			
			q_o			=> sipo_q,
			full_o		=> sipo_full
			);
			
			-- SIPO -- SB ->-> => SA
			sipo_d 		<= B_DAT_i;
			A_DAT_o 	<= sipo_q;
			sipo_sh_in 	<= B_ACK_i;
			sipo_clr 	<= sipo_full;
			A_ACK_o		<= sipo_full;
						
			process (clk_i)
			begin
				if (clk_i'event and clk_i = '1') then
					if(nRSt_i = '0') then
						--sipo_clr 	<= '0';
						sipo_sh_in 	<= '0';
						piso_ld 	<= '0';
						piso_sh_out	<= '0';
						B_CYC_o 	<= '0';
						B_STB_o 	<= '0';
						--A_ACK_o 	<= '0';
						A_STALL_o 	<= '0';
						CYC 		<= '0';
					else
						
						--sipo_clr 	<= '0';
						--sipo_sh_in 	<= '0';
						piso_ld 	<= '0';
						piso_sh_out	<= '0';
						B_CYC_o 	<= '0';
						B_STB_o 	<= '0';
						--A_ACK_o 	<= '0';
						A_STALL_o 	<= '0';
						
						CYC 		<= A_CYC_i;
						ld 			<= piso_ld;
						
						

						
						--piso_ld 
						if(A_STB_i = '1' AND piso_empty = '1') then
							piso_ld <= '1';
							--adr(A_ADR_i'left downto 0) <= A_ADR_i(A_ADR_i'left downto ld(g_dat_width_A/8-1)) & adr_zeros(ld(g_dat_width_A/8-1)-1 downto 0);
						end if;	
						
						
						
						--piso_sh_out
						if(B_STALL_i = '0' AND piso_empty = '0') then
							piso_sh_out <= '1';
							--adr <= adr + g_A_dat_width/8;
						end if;	
						
						-- CYC
						if(A_CYC_i = '1' OR piso_empty = '0') then
							B_CYC_o <= '1';
						end if;
						
						-- STB
						-- STALL						
						if(piso_empty = '0') then--falling edge
							B_STB_o <= '1';
							A_STALL_o <= '1';
						end if;	

						
						
						
						
						
					end if;	
				end if;
			end process;
				
		end GENERATE;

end architecture;